library IEEE;
use IEEE.std_logic_1164.all; -- import std_logic types
use IEEE.std_logic_arith.all; -- import add/sub of std_logic_vector
use IEEE.std_logic_unsigned.all;

use work.RISC_lib.all;

entity hazard_detect_unit is
	port ( id_ex_op1	:in data_word
						
				
		
		
		
		);
end hazard_detect_unit;

architecture behavioral of hazard_detect_unit is
begin
	process (id_ex_op1)
	begin
	
	end process;
end architecture behavioral;
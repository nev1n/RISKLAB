library IEEE;
use IEEE.std_logic_1164.all; -- import std_logic types
use IEEE.std_logic_arith.all; -- import add/sub of std_logic_vector
use IEEE.std_logic_unsigned.all;

use work.RISC_lib.all;

entity forward_unit is
	port (clk	:in std_logic
		);
end forward_unit;

architecture behavioral of forward_unit is
begin
	process (clk)
	begin
	
	end process;
end architecture behavioral;